
module uart_rx(

);

// receiver states /////////////////////////////////////////////////////////////
// localparam RESET = 0;
// localparam 


endmodule