module monitor_fpga(

);


endmodule