module monitor_fpga(
    input clk
);


endmodule