// uart.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module uart (
		input  wire        clk_clk,                        //                        clk.clk
		input  wire        reset_reset_n,                  //                      reset.reset_n
		input  wire        uart_0_external_connection_rxd, // uart_0_external_connection.rxd
		output wire        uart_0_external_connection_txd, //                           .txd
		output wire        uart_0_irq_irq,                 //                 uart_0_irq.irq
		input  wire [2:0]  uart_0_s1_address,              //                  uart_0_s1.address
		input  wire        uart_0_s1_begintransfer,        //                           .begintransfer
		input  wire        uart_0_s1_chipselect,           //                           .chipselect
		input  wire        uart_0_s1_read_n,               //                           .read_n
		input  wire        uart_0_s1_write_n,              //                           .write_n
		input  wire [15:0] uart_0_s1_writedata,            //                           .writedata
		output wire [15:0] uart_0_s1_readdata              //                           .readdata
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> uart_0:reset_n

	uart_uart_0 uart_0 (
		.clk           (clk_clk),                         //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset), //               reset.reset_n
		.address       (uart_0_s1_address),               //                  s1.address
		.begintransfer (uart_0_s1_begintransfer),         //                    .begintransfer
		.chipselect    (uart_0_s1_chipselect),            //                    .chipselect
		.read_n        (uart_0_s1_read_n),                //                    .read_n
		.write_n       (uart_0_s1_write_n),               //                    .write_n
		.writedata     (uart_0_s1_writedata),             //                    .writedata
		.readdata      (uart_0_s1_readdata),              //                    .readdata
		.rxd           (uart_0_external_connection_rxd),  // external_connection.export
		.txd           (uart_0_external_connection_txd),  //                    .export
		.irq           (uart_0_irq_irq)                   //                 irq.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
